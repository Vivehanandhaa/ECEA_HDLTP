`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 30.10.2022 02:17:21
// Design Name: 
// Module Name: exp_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module exp_tb;
reg A,B,C;
wire X;
exp uut (.A(A),.B(B),.C(C),.X(X));
initial begin
A=1'b0;B=1'b0;C=1'b0; #30
A=1'b0;B=1'b0;C=1'b1; #30
A=1'b0;B=1'b1;C=1'b0; #30
A=1'b0;B=1'b1;C=1'b1; #30
A=1'b1;B=1'b0;C=1'b0; #30
A=1'b1;B=1'b0;C=1'b1; #30
A=1'b1;B=1'b1;C=1'b0; #30
A=1'b1;B=1'b1;C=1'b1;
end
endmodule
